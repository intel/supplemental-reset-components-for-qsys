/*
 * Copyright (c) 2021 Intel Corporation
 *
 * SPDX-License-Identifier: MIT-0
 */

module sim_top ();

    test_sys_tb tb();
    sim_driver drvr();

endmodule
